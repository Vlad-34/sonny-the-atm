library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity sonny is
	
end sonny;

architecture structural of sonny is
begin
	
end structural;